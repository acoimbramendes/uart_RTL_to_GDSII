`include "uvm_macros.svh"
package uart_test_pkg;
	
	import uvm_pkg::*;
	
	`include "uart_transaction.sv"
	`include "drivers.sv"
	`include "monitors.sv"
	
endpackage: uart_test_pkg